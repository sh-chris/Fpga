
module niosIIsystem (
	clk_clk);	

	input		clk_clk;
endmodule
