// niosIIsystem.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module niosIIsystem (
		input  wire  clk_clk  // clk.clk
	);

	wire         nios2_core_debug_reset_request_reset;                      // nios2_core:debug_reset_request -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire  [31:0] nios2_core_data_master_readdata;                           // mm_interconnect_0:nios2_core_data_master_readdata -> nios2_core:d_readdata
	wire         nios2_core_data_master_waitrequest;                        // mm_interconnect_0:nios2_core_data_master_waitrequest -> nios2_core:d_waitrequest
	wire         nios2_core_data_master_debugaccess;                        // nios2_core:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_core_data_master_debugaccess
	wire  [13:0] nios2_core_data_master_address;                            // nios2_core:d_address -> mm_interconnect_0:nios2_core_data_master_address
	wire   [3:0] nios2_core_data_master_byteenable;                         // nios2_core:d_byteenable -> mm_interconnect_0:nios2_core_data_master_byteenable
	wire         nios2_core_data_master_read;                               // nios2_core:d_read -> mm_interconnect_0:nios2_core_data_master_read
	wire         nios2_core_data_master_readdatavalid;                      // mm_interconnect_0:nios2_core_data_master_readdatavalid -> nios2_core:d_readdatavalid
	wire         nios2_core_data_master_write;                              // nios2_core:d_write -> mm_interconnect_0:nios2_core_data_master_write
	wire  [31:0] nios2_core_data_master_writedata;                          // nios2_core:d_writedata -> mm_interconnect_0:nios2_core_data_master_writedata
	wire  [31:0] nios2_core_instruction_master_readdata;                    // mm_interconnect_0:nios2_core_instruction_master_readdata -> nios2_core:i_readdata
	wire         nios2_core_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_core_instruction_master_waitrequest -> nios2_core:i_waitrequest
	wire  [12:0] nios2_core_instruction_master_address;                     // nios2_core:i_address -> mm_interconnect_0:nios2_core_instruction_master_address
	wire         nios2_core_instruction_master_read;                        // nios2_core:i_read -> mm_interconnect_0:nios2_core_instruction_master_read
	wire         nios2_core_instruction_master_readdatavalid;               // mm_interconnect_0:nios2_core_instruction_master_readdatavalid -> nios2_core:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:Jtag_uart_avalon_jtag_slave_chipselect -> Jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // Jtag_uart:av_readdata -> mm_interconnect_0:Jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // Jtag_uart:av_waitrequest -> mm_interconnect_0:Jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:Jtag_uart_avalon_jtag_slave_address -> Jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:Jtag_uart_avalon_jtag_slave_read -> Jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:Jtag_uart_avalon_jtag_slave_write -> Jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:Jtag_uart_avalon_jtag_slave_writedata -> Jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_systemid_control_slave_readdata;         // systemID:readdata -> mm_interconnect_0:systemID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_systemid_control_slave_address;          // mm_interconnect_0:systemID_control_slave_address -> systemID:address
	wire  [31:0] mm_interconnect_0_nios2_core_debug_mem_slave_readdata;     // nios2_core:debug_mem_slave_readdata -> mm_interconnect_0:nios2_core_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_core_debug_mem_slave_waitrequest;  // nios2_core:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_core_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_core_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_core_debug_mem_slave_debugaccess -> nios2_core:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_core_debug_mem_slave_address;      // mm_interconnect_0:nios2_core_debug_mem_slave_address -> nios2_core:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_core_debug_mem_slave_read;         // mm_interconnect_0:nios2_core_debug_mem_slave_read -> nios2_core:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_core_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_core_debug_mem_slave_byteenable -> nios2_core:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_core_debug_mem_slave_write;        // mm_interconnect_0:nios2_core_debug_mem_slave_write -> nios2_core:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_core_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_core_debug_mem_slave_writedata -> nios2_core:debug_mem_slave_writedata
	wire         mm_interconnect_0_sram_s1_chipselect;                      // mm_interconnect_0:SRAM_s1_chipselect -> SRAM:chipselect
	wire  [31:0] mm_interconnect_0_sram_s1_readdata;                        // SRAM:readdata -> mm_interconnect_0:SRAM_s1_readdata
	wire   [9:0] mm_interconnect_0_sram_s1_address;                         // mm_interconnect_0:SRAM_s1_address -> SRAM:address
	wire   [3:0] mm_interconnect_0_sram_s1_byteenable;                      // mm_interconnect_0:SRAM_s1_byteenable -> SRAM:byteenable
	wire         mm_interconnect_0_sram_s1_write;                           // mm_interconnect_0:SRAM_s1_write -> SRAM:write
	wire  [31:0] mm_interconnect_0_sram_s1_writedata;                       // mm_interconnect_0:SRAM_s1_writedata -> SRAM:writedata
	wire         mm_interconnect_0_sram_s1_clken;                           // mm_interconnect_0:SRAM_s1_clken -> SRAM:clken
	wire         irq_mapper_receiver0_irq;                                  // Jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_core_irq_irq;                                        // irq_mapper:sender_irq -> nios2_core:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [Jtag_uart:rst_n, irq_mapper:reset, mm_interconnect_0:nios2_core_reset_reset_bridge_in_reset_reset, nios2_core:reset_n, rst_translator:in_reset, systemID:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [nios2_core:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [SRAM:reset, mm_interconnect_0:SRAM_reset1_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> SRAM:reset_req

	niosIIsystem_Jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	niosIIsystem_SRAM sram (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_sram_s1_address),      //     s1.address
		.clken      (mm_interconnect_0_sram_s1_clken),        //       .clken
		.chipselect (mm_interconnect_0_sram_s1_chipselect),   //       .chipselect
		.write      (mm_interconnect_0_sram_s1_write),        //       .write
		.readdata   (mm_interconnect_0_sram_s1_readdata),     //       .readdata
		.writedata  (mm_interconnect_0_sram_s1_writedata),    //       .writedata
		.byteenable (mm_interconnect_0_sram_s1_byteenable),   //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)  //       .reset_req
	);

	niosIIsystem_nios2_core nios2_core (
		.clk                                 (clk_clk),                                                  //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                          //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                       //                          .reset_req
		.d_address                           (nios2_core_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_core_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_core_data_master_read),                              //                          .read
		.d_readdata                          (nios2_core_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_core_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_core_data_master_write),                             //                          .write
		.d_writedata                         (nios2_core_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_core_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_core_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_core_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_core_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_core_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_core_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_core_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_core_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_core_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_core_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_core_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_core_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_core_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_core_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_core_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_core_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_core_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	niosIIsystem_systemID systemid (
		.clock    (clk_clk),                                           //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_systemid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_systemid_control_slave_address)   //              .address
	);

	niosIIsystem_mm_interconnect_0 mm_interconnect_0 (
		.main_clock_clk_clk                           (clk_clk),                                                   //                         main_clock_clk.clk
		.nios2_core_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // nios2_core_reset_reset_bridge_in_reset.reset
		.SRAM_reset1_reset_bridge_in_reset_reset      (rst_controller_001_reset_out_reset),                        //      SRAM_reset1_reset_bridge_in_reset.reset
		.nios2_core_data_master_address               (nios2_core_data_master_address),                            //                 nios2_core_data_master.address
		.nios2_core_data_master_waitrequest           (nios2_core_data_master_waitrequest),                        //                                       .waitrequest
		.nios2_core_data_master_byteenable            (nios2_core_data_master_byteenable),                         //                                       .byteenable
		.nios2_core_data_master_read                  (nios2_core_data_master_read),                               //                                       .read
		.nios2_core_data_master_readdata              (nios2_core_data_master_readdata),                           //                                       .readdata
		.nios2_core_data_master_readdatavalid         (nios2_core_data_master_readdatavalid),                      //                                       .readdatavalid
		.nios2_core_data_master_write                 (nios2_core_data_master_write),                              //                                       .write
		.nios2_core_data_master_writedata             (nios2_core_data_master_writedata),                          //                                       .writedata
		.nios2_core_data_master_debugaccess           (nios2_core_data_master_debugaccess),                        //                                       .debugaccess
		.nios2_core_instruction_master_address        (nios2_core_instruction_master_address),                     //          nios2_core_instruction_master.address
		.nios2_core_instruction_master_waitrequest    (nios2_core_instruction_master_waitrequest),                 //                                       .waitrequest
		.nios2_core_instruction_master_read           (nios2_core_instruction_master_read),                        //                                       .read
		.nios2_core_instruction_master_readdata       (nios2_core_instruction_master_readdata),                    //                                       .readdata
		.nios2_core_instruction_master_readdatavalid  (nios2_core_instruction_master_readdatavalid),               //                                       .readdatavalid
		.Jtag_uart_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //            Jtag_uart_avalon_jtag_slave.address
		.Jtag_uart_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                       .write
		.Jtag_uart_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                       .read
		.Jtag_uart_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                       .readdata
		.Jtag_uart_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                       .writedata
		.Jtag_uart_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                       .waitrequest
		.Jtag_uart_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                       .chipselect
		.nios2_core_debug_mem_slave_address           (mm_interconnect_0_nios2_core_debug_mem_slave_address),      //             nios2_core_debug_mem_slave.address
		.nios2_core_debug_mem_slave_write             (mm_interconnect_0_nios2_core_debug_mem_slave_write),        //                                       .write
		.nios2_core_debug_mem_slave_read              (mm_interconnect_0_nios2_core_debug_mem_slave_read),         //                                       .read
		.nios2_core_debug_mem_slave_readdata          (mm_interconnect_0_nios2_core_debug_mem_slave_readdata),     //                                       .readdata
		.nios2_core_debug_mem_slave_writedata         (mm_interconnect_0_nios2_core_debug_mem_slave_writedata),    //                                       .writedata
		.nios2_core_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_core_debug_mem_slave_byteenable),   //                                       .byteenable
		.nios2_core_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_core_debug_mem_slave_waitrequest),  //                                       .waitrequest
		.nios2_core_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_core_debug_mem_slave_debugaccess),  //                                       .debugaccess
		.SRAM_s1_address                              (mm_interconnect_0_sram_s1_address),                         //                                SRAM_s1.address
		.SRAM_s1_write                                (mm_interconnect_0_sram_s1_write),                           //                                       .write
		.SRAM_s1_readdata                             (mm_interconnect_0_sram_s1_readdata),                        //                                       .readdata
		.SRAM_s1_writedata                            (mm_interconnect_0_sram_s1_writedata),                       //                                       .writedata
		.SRAM_s1_byteenable                           (mm_interconnect_0_sram_s1_byteenable),                      //                                       .byteenable
		.SRAM_s1_chipselect                           (mm_interconnect_0_sram_s1_chipselect),                      //                                       .chipselect
		.SRAM_s1_clken                                (mm_interconnect_0_sram_s1_clken),                           //                                       .clken
		.systemID_control_slave_address               (mm_interconnect_0_systemid_control_slave_address),          //                 systemID_control_slave.address
		.systemID_control_slave_readdata              (mm_interconnect_0_systemid_control_slave_readdata)          //                                       .readdata
	);

	niosIIsystem_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_core_irq_irq)              //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_core_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (nios2_core_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),       // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),   //          .reset_req
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_core_debug_reset_request_reset),   // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
